
module top_tb;

endmodule : top_tb
